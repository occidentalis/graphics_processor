module rasterizer_unit (
	input logic [47:0] p1, p2, p3,
	input logic [15:0] pixel_x, pixel_y,
	
);