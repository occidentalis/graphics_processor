module shader_unit (
    input logic clk, start,
    input logic [31:0] p1[3], p2[3], p3[3], // in NDC coordinates
    output logic [3:0] color,
    output logic done
);



endmodule